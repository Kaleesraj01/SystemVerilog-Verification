interface intf;
  logic [3:0]din;
  logic clk , rst ;
  logic [3:0]q ;
 
endinterface 
