 interface intf;
 
  (
     logic clk,
      logic rst_n,
     logic [3:0] count );
endinterface 
